module DE10 (
	input CLOCK_50,
	input [3:0] KEY,
	output [9:0] LEDR
);

	
endmodule